module test (
    input clk,
    input rst


);
  assign clk = rst;
endmodule

